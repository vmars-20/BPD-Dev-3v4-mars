--------------------------------------------------------------------------------
-- File: CustomWrapper_bpd_forge.vhd
-- Author: Moku Instrument Forge Team
-- Date: 2025-11-05
-- Version: 3.0 (Forge 3-layer architecture)
--
-- Description:
--   CustomWrapper architecture for Basic Probe Driver using Forge 3-layer pattern.
--   Implements FORGE_READY control scheme (CR0[31:29]) for safe MCC integration.
--
-- Entity: CustomWrapper (defined in CustomWrapper_test_stub.vhd)
--
-- FORGE Control Scheme (CR0[31:29]):
--   CR0[31] = forge_ready  - Set by MCC loader after deployment
--   CR0[30] = user_enable  - User control (GUI toggle)
--   CR0[29] = clk_enable   - Clock gating control
--   loader_done            - BRAM loader completion (tied to '1' for now)
--
-- Register Mapping:
--   CR0[31:29] → FORGE control bits (3-bit handshaking)
--   CR1-CR11   → Application registers (11 registers)
--
-- Architecture:
--   Layer 1: (MCC_TOP_forge_loader.vhd - future)
--   Layer 2: BPD_forge_shim.vhd (register mapping)
--   Layer 3: BPD_forge_main.vhd (FSM logic)
--
-- Platform: Moku:Go
-- Clock Frequency: 125 MHz
--
-- References:
--   - forge_common_pkg.vhd (FORGE_READY control scheme)
--   - BPD_forge_shim.vhd (shim layer)
--   - BPD_forge_main.vhd (main logic)
--   - external_Example/DS1140_polo_shim.vhd (pattern reference)
--------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

architecture bpd_forge of CustomWrapper is

    ----------------------------------------------------------------------------
    -- FORGE Control Signals (extracted from CR0[31:29])
    ----------------------------------------------------------------------------
    signal forge_ready  : std_logic;
    signal user_enable  : std_logic;
    signal clk_enable   : std_logic;
    signal loader_done  : std_logic;

begin

    ----------------------------------------------------------------------------
    -- Extract FORGE Control Bits from Control0
    --
    -- CR0[31] = forge_ready  (set by loader after deployment)
    -- CR0[30] = user_enable  (user control)
    -- CR0[29] = clk_enable   (clock gating)
    ----------------------------------------------------------------------------
    forge_ready <= Control0(31);
    user_enable <= Control0(30);
    clk_enable  <= Control0(29);

    ----------------------------------------------------------------------------
    -- BRAM Loader Done Signal
    --
    -- TODO: Connect to actual BRAM loader when implemented
    -- For now, tie to '1' (no BRAM loading required)
    ----------------------------------------------------------------------------
    loader_done <= '1';

    ----------------------------------------------------------------------------
    -- Instantiate BPD Forge Shim (Layer 2)
    --
    -- The shim layer:
    --   1. Receives FORGE control signals
    --   2. Maps app_reg_1..app_reg_11 to friendly names
    --   3. Computes global_enable via combine_forge_ready()
    --   4. Instantiates BPD_forge_main (Layer 3)
    ----------------------------------------------------------------------------
    BPD_SHIM_INST: entity WORK.BPD_forge_shim
        port map (
            -- Clock and Reset
            Clk   => Clk,
            Reset => Reset,

            -- FORGE Control (3-bit handshaking scheme)
            forge_ready  => forge_ready,
            user_enable  => user_enable,
            clk_enable   => clk_enable,
            loader_done  => loader_done,

            -- Application Registers (CR1-CR11)
            app_reg_1  => Control1,
            app_reg_2  => Control2,
            app_reg_3  => Control3,
            app_reg_4  => Control4,
            app_reg_5  => Control5,
            app_reg_6  => Control6,
            app_reg_7  => Control7,
            app_reg_8  => Control8,
            app_reg_9  => Control9,
            app_reg_10 => Control10,
            app_reg_11 => Control11,

            -- BRAM Interface (reserved for future use)
            bram_addr => (others => '0'),
            bram_data => (others => '0'),
            bram_we   => '0',

            -- MCC I/O (FORGE Standard: 2 inputs, 3 outputs)
            -- InputC reserved for BRAM loader (future)
            -- OutputC driven by SHIM hierarchical encoder
            InputA  => InputA,
            InputB  => InputB,
            OutputA => OutputA,
            OutputB => OutputB,
            OutputC => OutputC
        );

end architecture bpd_forge;

--------------------------------------------------------------------------------
-- Usage Instructions
--------------------------------------------------------------------------------
--
-- 1. FORGE Control Initialization Sequence:
--
--    a) Power-on: Control0 = 0x00000000
--       → forge_ready=0, user_enable=0, clk_enable=0
--       → Module disabled (safe default)
--
--    b) MCC loader sets Control0[31] = 1
--       → forge_ready=1 (deployment complete)
--
--    c) User enables module via GUI: Control0[30] = 1
--       → user_enable=1
--
--    d) User enables clock: Control0[29] = 1
--       → clk_enable=1
--
--    e) Module operates: global_enable = forge_ready AND user_enable AND clk_enable AND loader_done
--
-- 2. Application Register Mapping (CR1-CR11):
--
--    CR1[3:0]   : Lifecycle control (arm_enable, ext_trigger_in, auto_rearm, fault_clear)
--    CR2[15:0]  : Trigger output voltage (mV)
--    CR3[15:0]  : Trigger pulse duration (ns)
--    CR4[15:0]  : Intensity output voltage (mV)
--    CR5[15:0]  : Intensity pulse duration (ns)
--    CR6[15:0]  : Trigger wait timeout (s)
--    CR7[23:0]  : Cooldown interval (μs)
--    CR8[1:0]   : Monitor control (enable, expect_negative)
--    CR9[15:0]  : Monitor threshold voltage (mV)
--    CR10[31:0] : Monitor window start delay (ns)
--    CR11[31:0] : Monitor window duration (ns)
--
-- 3. MCC I/O Mapping:
--
--    InputA  → probe_monitor_feedback (ADC, ±5V)
--    InputB  → (unused)
--    OutputA → Trigger output (DAC, ±5V)
--    OutputB → Intensity output (DAC, ±5V)
--    OutputC → (reserved)
--    OutputD → Hierarchical voltage encoding (FSM state + app status, debugging)
--
-- 4. Hierarchical Voltage Encoding (OutputD):
--
--    NEW (Handoff 6): OutputD driven by SHIM layer with hierarchical encoder
--    - Encodes 14 bits: 6-bit FSM state + 8-bit app status
--    - Major transitions: 200 digital units per state (human-readable on scope)
--    - Status information: Fine-grained offset (machine-decodable)
--    - Fault detection: Negative voltage (status[7] = fault flag)
--    - Replaces: fsm_observer.vhd LUT-based pattern
--    - Benefits: Zero LUTs, 14-bit density, single bitstream dev/prod
--
--    Reference: Obsidian/Project/Handoffs/2025-11-07-handoff-6-hierarchical-voltage-encoding.md
--
--------------------------------------------------------------------------------
